LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.std_logic_arith.ALL;

ENTITY datapath IS
	GENERIC (
		DATA_WIDTH : INTEGER := 16;
		ADDR_WIDTH : INTEGER := 4
	);
	PORT (
		rst : IN STD_LOGIC;
		clk : IN STD_LOGIC;
		imm : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		data_in_mux2 : IN STD_LOGIC_VECTOR(DATA_WIDTH - 1 DOWNTO 0);
		RFs : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		ALUs : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		ALUz : OUT STD_LOGIC;
		ALUeq : OUT STD_LOGIC;
		ALUgt : OUT STD_LOGIC;

		RFwa : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		RFwe : IN STD_LOGIC;
		OPr1a : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		OPr1e : IN STD_LOGIC;
		OPr2a : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		OPr2e : IN STD_LOGIC;

		add_out : OUT STD_LOGIC_VECTOR(DATA_WIDTH - 1 DOWNTO 0);
		data_out : OUT STD_LOGIC_VECTOR(DATA_WIDTH - 1 DOWNTO 0)
	);
END datapath;

ARCHITECTURE struct OF datapath IS
	COMPONENT alu
		PORT (
			OPr1 : IN STD_LOGIC_VECTOR(DATA_WIDTH - 1 DOWNTO 0);
			OPr2 : IN STD_LOGIC_VECTOR(DATA_WIDTH - 1 DOWNTO 0);
			ALUs : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			ALUz : OUT STD_LOGIC;
			ALUeq : OUT STD_LOGIC;
			ALUgt : OUT STD_LOGIC;
			ALUr : OUT STD_LOGIC_VECTOR(DATA_WIDTH - 1 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT mux4to1
		GENERIC (DATA_WIDTH : INTEGER := 16);
		PORT (
			data_in_mux0, data_in_mux1, data_in_mux2, data_in_mux3 : IN STD_LOGIC_VECTOR (DATA_WIDTH - 1 DOWNTO 0);
			SEL : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
			Z : OUT STD_LOGIC_VECTOR (DATA_WIDTH - 1 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT register_file
		GENERIC (
			DATA_WIDTH : INTEGER := 16;
			ADDR_WIDTH : INTEGER := 4
		);
		PORT (
			reset : IN STD_LOGIC;
			clk : IN STD_LOGIC;
			RFin : IN STD_LOGIC_VECTOR (DATA_WIDTH - 1 DOWNTO 0);
			RFwa : IN STD_LOGIC_VECTOR (ADDR_WIDTH - 1 DOWNTO 0);
			RFwe : IN STD_LOGIC;
			OPr1a : IN STD_LOGIC_VECTOR (ADDR_WIDTH - 1 DOWNTO 0);
			OPr1e : IN STD_LOGIC;
			OPr2a : IN STD_LOGIC_VECTOR (ADDR_WIDTH - 1 DOWNTO 0);
			OPr2e : IN STD_LOGIC;
			OPr1 : OUT STD_LOGIC_VECTOR (DATA_WIDTH - 1 DOWNTO 0);
			OPr2 : OUT STD_LOGIC_VECTOR (DATA_WIDTH - 1 DOWNTO 0));
	END COMPONENT;
	SIGNAL ALUr : STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL RFin : STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL data_in_mux3 : STD_LOGIC_VECTOR(15 DOWNTO 0) := x"0000";

	SIGNAL o1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL o2 : STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL data_in_mux1 : STD_LOGIC_VECTOR(15 DOWNTO 0);

BEGIN
	data_in_mux1 <= x"00" & imm;

	mux : mux4to1
	PORT MAP(ALUr, data_in_mux1, data_in_mux2, data_in_mux3, RFs, RFin);

	rf_u : register_file
	PORT MAP(rst, clk, RFin, RFwa, RFwe, OPr1a, OPr1e, OPr2a, OPr2e, o1, o2);

	alu_u : ALU
	PORT MAP(o1, o2, ALUs, ALUz, ALUeq, ALUgt, ALUr);
	add_out <= o2;
	data_out <= o1;

END struct;
